module not_op (x,f);
input x;
output f;
assign f=!x;
endmodule
